library verilog;
use verilog.vl_types.all;
entity AD_ctr_vlg_vec_tst is
end AD_ctr_vlg_vec_tst;
