library verilog;
use verilog.vl_types.all;
entity trigger_sec_vlg_vec_tst is
end trigger_sec_vlg_vec_tst;
