library verilog;
use verilog.vl_types.all;
entity measuring_vlg_vec_tst is
end measuring_vlg_vec_tst;
