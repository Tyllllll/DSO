library verilog;
use verilog.vl_types.all;
entity clk_generate_vlg_vec_tst is
end clk_generate_vlg_vec_tst;
