library verilog;
use verilog.vl_types.all;
entity measuring_vlg_sample_tst is
    port(
        clk             : in     vl_logic;
        data            : in     vl_logic_vector(9 downto 0);
        hscan_switch    : in     vl_logic;
        reset           : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end measuring_vlg_sample_tst;
